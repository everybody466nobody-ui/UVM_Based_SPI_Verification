interface spi_slave_if (input bit sck);
    
  
    logic mosi;
    logic miso;
    
    

endinterface

